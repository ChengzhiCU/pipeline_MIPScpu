module pipe_rom(reset,PC,enable,Instruction);
input reset,enable;
input [31:0] PC;
output wire [31:0] Instruction;
reg [31:0] Instruct;
assign Instruction = enable? Instruct:32'b0;
always@(*) 
 begin
	if(~reset) Instruct<=32'b0;
	else 
	 begin
		case(PC[30:2])
		/*
		0: Instruct <= 32'b001000_00000_10000_0000000000111011;  //addi $s0,$0,59
		1: Instruct <= 32'b001000_00000_10001_0000000001001011;  //addi $s1,$0,75
		2: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		3: Instruct <= 32'b000100_00000_10010_0000000000000111; //compare: beq $0,$s2,result
		4: Instruct <= 32'b000001_10010_00000_0000000000000011; //bltz $s2,neg
		5: Instruct <= 32'b000000_10000_10001_10000_00000_100010; //pos: sub $s0,$s0,$s1
		6: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		7: Instruct <= 32'b000010_00000000000000000000000011;    // j compare
		8: Instruct <= 32'b000000_10001_10000_10001_00000_100010; //neg: sub $s1,$s1,$s0
		9: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		10: Instruct <= 32'b000010_00000000000000000000000011;    // j compare
		11: Instruct <= 32'b101011_00100_10000_0000000000011000;  // result: sw $s0,00x0018($a0)
		*/
		
		
		0: Instruct <= 32'b000010_00000000000000000000000011; //j Normal
		1: Instruct <= 32'b000010_00000000000000000001101011; //j Interrupt
		2: Instruct <= 32'b000010_00000000000000000001101010;    //j Exit
		3: Instruct <= 32'b001111_00000_00100_1000000000000000;  //lui $a0,0x80000000
		4: Instruct <= 32'b001111_00000_00010_0000000000000000;  //lui $v0,0
		5: Instruct <= 32'b001111_00000_00011_0000000000000000;  //lui $v0,0
		6: Instruct <= 32'b000000_00000_00000_01000_00000_100000;//add $t0,$0,$0
		8: Instruct <= 32'b000000_00000_00000_01001_00000_100000;//add $t1,$0,$0
		7: Instruct <= 32'b001000_00000_00010_0000000000000010;  //addi $v0,$0,0x0002
		9: Instruct <= 32'b001000_00000_00011_0000000000001010;  //addi $v1,$0,0x000a
		
		10: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		
		11: Instruct <= 32'b100011_00100_01000_0000000000100000;   //loop1: lw $t0,0x0020($a0)
		
		15: Instruct <= 32'b000100_01000_00011_0000000000000101;  //beq $t0,$v1,break1
		
		20: Instruct <= 32'b000010_00000000000000000000001011;    // j loop1
		
		26: Instruct <= 32'b100011_00100_01001_0000000000011100;  //break1: lw $t1,0x001c($a0)
		
		31: Instruct = 32'b001000_00000_00010_0000000000000000;  //addi $v0,$0,0x0
		
		36: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		37: Instruct <= 32'b000000_00000_01001_10000_00000_100000; //add $s0,$0,$t1
		38: Instruct <= 32'b001000_00000_00010_0000000000000010;  //addi $v0,$0,0x0002
		
		39: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		
		40: Instruct <= 32'b100011_00100_01000_0000000000100000;   //loop2: lw $t0,0x0020($a0)
		45: Instruct <= 32'b000100_01000_00011_0000000000000101;  //beq $t0,$v1,break2
		50: Instruct <= 32'b000010_00000000000000000000101000;    // j loop2 
		56: Instruct <= 32'b100011_00100_01011_0000000000011100;  //break2: lw $t3,0x001c($a0)
		61: Instruct <= 32'b001000_00000_00010_0000000000000000;  //addi $v0,$0,0x0
		66: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		67: Instruct <= 32'b000000_00000_01011_10001_00000_100000; //add $s1,$0,$t3
		
		68: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		69: Instruct <= 32'b000100_00000_10010_0000000000000111; //compare: beq $0,$s2,result
		70: Instruct <= 32'b000001_10010_00000_0000000000000011; //bltz $s2,neg
		71: Instruct <= 32'b000000_10000_10001_10000_00000_100010; //pos: sub $s0,$s0,$s1
		72: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		73: Instruct <= 32'b000010_00000000000000000001000101;    // j compare
		74: Instruct <= 32'b000000_10001_10000_10001_00000_100010; //neg: sub $s1,$s1,$s0
		75: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		76: Instruct <= 32'b000010_00000000000000000001000101;    // j compare
		77: Instruct <= 32'b101011_00100_10000_0000000000011000;  // result: sw $s0,00x0018($a0)
		
		82: Instruct <= 32'b001000_00000_00010_0000000000000001;  //addi $v0,$0,0x0001
		83: Instruct <= 32'b001000_00000_00011_0000000000000101;  //addi $v1,$0,0x0005
		84: Instruct <= 32'b101011_00100_00010_0000000000100000;  //sw $v0,0x0020($a0)
		85: Instruct <= 32'b100011_00100_01010_0000000000100000;   //loop3: lw $t2,0x0020($a0)
		86: Instruct <= 32'b000100_01010_00011_0000000000000101;  //beq $t2,$v1,break3
		91: Instruct <= 32'b000010_00000000000000000001010101;    // j loop3
		97: Instruct <= 32'b001000_00000_00010_0000000000000000;  //break3:addi $v0,$0,0x0000
		102: Instruct <= 32'b101011_00100_00010_0000000000100000;  //sw $v0,0x0020($a0)
		103: Instruct <= 32'b001111_00000_00100_0100000000000000;  //lui $a0,0x40000000
		108: Instruct <= 32'b101011_00100_10000_0000000000001100;  //sw $s0,0x000c($a0) 
		
		/*
		47: Instruct <= 32'b001000_00000_00010_0000000000000001;  //addi $v0,$0,0x0001
		48: Instruct <= 32'b101011_00000_00010_0000000000000000;  //sw $v0,0x0000($0)
		49: Instruct <= 32'b001000_00000_00010_0000000001001111;  //addi $v0,$0,0x004f
		50: Instruct <= 32'b101011_00000_00010_0000000000000100;  //sw $v0,0x0004($0)
		51: Instruct <= 32'b001000_00000_00010_0000000000010010;  //addi $v0,$0,0x0012
		52: Instruct <= 32'b101011_00000_00010_0000000000001000;  //sw $v0,0x0008($0)
		53: Instruct <= 32'b001000_00000_00010_0000000000000110;  //addi $v0,$0,0x0006
		54: Instruct <= 32'b101011_00000_00010_0000000000001100;  //sw $v0,0x000c($0)
		55: Instruct <= 32'b001000_00000_00010_0000000001001100;  //addi $v0,$0,0x004c
		56: Instruct <= 32'b101011_00000_00010_0000000000010000;  //sw $v0,0x0010($0)
		57: Instruct <= 32'b001000_00000_00010_0000000000100100;  //addi $v0,$0,0x0024
		58: Instruct <= 32'b101011_00000_00010_0000000000010100;  //sw $v0,0x0014($0)
		59: Instruct <= 32'b001000_00000_00010_0000000000100000;  //addi $v0,$0,0x0020
		60: Instruct <= 32'b101011_00000_00010_0000000000011000;  //sw $v0,0x0018($0)
		61: Instruct <= 32'b001000_00000_00010_0000000000001111;  //addi $v0,$0,0x000f
		62: Instruct <= 32'b101011_00000_00010_0000000000011100;  //sw $v0,0x001c($0)
		63: Instruct <= 32'b001000_00000_00010_0000000000000000;  //addi $v0,$0,0x0000
		64: Instruct <= 32'b101011_00000_00010_0000000000100000;  //sw $v0,0x0020($0)
		65: Instruct <= 32'b001000_00000_00010_0000000000000100;  //addi $v0,$0,0x0004
		66: Instruct <= 32'b101011_00000_00010_0000000000100100;  //sw $v0,0x0024($0)
		67: Instruct <= 32'b001000_00000_00010_0000000000001000;  //addi $v0,$0,0x0008
		68: Instruct <= 32'b101011_00000_00010_0000000000101000;  //sw $v0,0x0028($0)
		69: Instruct <= 32'b001000_00000_00010_0000000001100000;  //addi $v0,$0,0x0060
		70: Instruct <= 32'b101011_00000_00010_0000000000101100;  //sw $v0,0x002c($0)
		71: Instruct <= 32'b001000_00000_00010_0000000000110001;  //addi $v0,$0,0x0031
		72: Instruct <= 32'b101011_00000_00010_0000000000110000;  //sw $v0,0x0030($0)
		73: Instruct <= 32'b001000_00000_00010_0000000001000010;  //addi $v0,$0,0x0042
		74: Instruct <= 32'b101011_00000_00010_0000000000110100;  //sw $v0,0x0034($0)
		75: Instruct <= 32'b001000_00000_00010_0000000000110000;  //addi $v0,$0,0x0030
		76: Instruct <= 32'b101011_00000_00010_0000000000111000;  //sw $v0,0x0038($0)
		77: Instruct <= 32'b001000_00000_00010_0000000000111000;  //addi $v0,$0,0x0038
		78: Instruct <= 32'b101011_00000_00010_0000000000111100;  //sw $v0,0x003c($0)
		79: Instruct <= 32'b000000_00000_00000_00010_00000_100000;//add $v0,$0,$0
		80: Instruct <= 32'b101011_00100_00010_0000000000001000;  //sw,$v0,0x0008($a0)
		81: Instruct <= 32'b001111_00000_00010_1111111111111111;  //lui $v0,0xffff
		82: Instruct <= 32'b001001_00010_00010_1111111111111111;  //addiu $v0,$v0,0xffff
		83: Instruct <= 32'b101011_00100_00010_0000000000000100;  //sw,$v0,0x0004($a0)
		84: Instruct <= 32'b001000_00000_00010_1111111100000000;  //addi $v0,$0,0xff00
		85: Instruct <= 32'b0;  //nop
		86: Instruct <= 32'b101011_00100_00010_0000000000000000;  //sw $v0,0x0000($a0)
		87: Instruct <= 32'b001100_01001_10000_0000000000001111;  //andi $s0,$t1,0x000f
		88: Instruct <= 32'b001100_01001_10001_0000000011110000;  //andi $s1,$t1,0x00f0
		89: Instruct <= 32'b000000_00000_10001_10001_00010_000010;//srl $s1,$s1,2
		90: Instruct <= 32'b001100_01011_10010_0000000000001111;  //andi $s0,$t1,0x000f
		91: Instruct <= 32'b001100_01011_10011_0000000011110000;  //andi $s1,$t1,0x00f0
		92: Instruct <= 32'b000000_00000_10011_10011_00010_000010;//srl $s1,$s1,2
		93: Instruct <= 32'b000000_00000_10000_10000_00010_000000;//sll $s0,$s0,2
		94: Instruct <= 32'b000000_00000_10010_10010_00010_000000;//sll $s2,$s2,2
		95: Instruct <= 32'b100011_10000_10000_0000000000000000;  //lw $s0,0x0000($s0)
		96: Instruct <= 32'b100011_10001_10001_0000000000000000;  //lw $s1,0x0000($s1)
		97: Instruct <= 32'b100011_10010_10010_0000000000000000;  //lw $s2,0x0000($s2)
		98: Instruct <= 32'b100011_10011_10011_0000000000000000;  //lw $s3,0x0000($s3)
		99: Instruct <= 32'b001000_00000_11000_0000000100000000;  //addi $t8,$0,0x0100
		100: Instruct <= 32'b001000_00000_10100_0000000100000000;  //addi $s4,$0,0x0100
		101: Instruct <= 32'b001000_00000_10101_0000001000000000;  //addi $s5,$0,0x0200
		102: Instruct <= 32'b001000_00000_10110_0000010000000000;  //addi $s6,$0,0x0400
		103: Instruct <= 32'b001000_00000_10111_0000100000000000;  //addi $s7,$0,0x0800
		104: Instruct <= 32'b001000_00000_00010_0000000000000011;  //addi $v0,$0,0x0003
		105: Instruct <= 32'b101011_00100_00010_0000000000001000;  //sw $v0,0x0008($a0)
		106: Instruct <= 32'b0;    //Exit: j Exit
		107: Instruct <= 32'b001000_00000_00011_0000000000000001;  //Interrupt: addi $v1,$0,0x0001
		108: Instruct <= 32'b101011_00100_00011_0000000000001000;  //sw $v1,0x0008($a0)
		109: Instruct <= 32'b000100_11000_10100_0000000000000011;  //beq $t8,$s4,one
		110: Instruct <= 32'b000100_11000_10101_0000000000001000;  //beq $t8,$s5,two
		111: Instruct <= 32'b000100_11000_10110_0000000000001101;  //beq $t8,$s6,three
		112: Instruct <= 32'b000100_11000_10111_0000000000010010;  //beq $t8,$s7,four
		113: Instruct <= 32'b000000_11000_10000_00010_00000_100000;//one: add $v0,$t8,$s0
		114: Instruct <= 32'b101011_00100_00010_0000000000010100;  //sw $v0,0x0014($a0)
		115: Instruct <= 32'b001000_00000_11000_0000001000000000;  //addi $t8,$0,0x0200
		116: Instruct <= 32'b001000_00000_00011_0000000000000011;  //addi $v1,$0,0x0003
		117: Instruct <= 32'b101011_00100_00011_0000000000001000;  //sw $v1,0x0008($a0)
		118: Instruct <= 32'b000000_11010_00000_00000_00000_001000;//jr $26
		119: Instruct <= 32'b000000_11000_10001_00010_00000_100000;//two: add $v0,$t8,$s1
		120: Instruct <= 32'b101011_00100_00010_0000000000010100;  //sw $v0,0x0014($a0)
		121: Instruct <= 32'b001000_00000_11000_0000010000000000;  //addi $t8,$0,0x0400
		122: Instruct <= 32'b001000_00000_00011_0000000000000011;  //addi $v1,$0,0x0003
		123: Instruct <= 32'b101011_00100_00011_0000000000001000;  //sw $v1,0x0008($a0)
		124: Instruct <= 32'b000000_11010_00000_00000_00000_001000;//jr $26
		125: Instruct <= 32'b000000_11000_10010_00010_00000_100000;//three: add $v0,$t8,$s2
		126: Instruct <= 32'b101011_00100_00010_0000000000010100;  //sw $v0,0x0014($a0)
		127: Instruct <= 32'b001000_00000_11000_0000100000000000;  //addi $t8,$0,0x0800
		128: Instruct <= 32'b001000_00000_00011_0000000000000011;  //addi $v1,$0,0x0003
		129: Instruct <= 32'b101011_00100_00011_0000000000001000;  //sw $v1,0x0008($a0)
		130: Instruct <= 32'b000000_11010_00000_00000_00000_001000;//jr $26
		131: Instruct <= 32'b000000_11000_10011_00010_00000_100000;//one: add $v0,$t8,$s3
		132: Instruct <= 32'b101011_00100_00010_0000000000010100;  //sw $v0,0x0014($a0)
		133: Instruct <= 32'b001000_00000_11000_0000000100000000;  //addi $t8,$0,0x0100
		134: Instruct <= 32'b001000_00000_00011_0000000000000011;  //addi $v1,$0,0x0003
		135: Instruct <= 32'b101011_00100_00011_0000000000001000;  //sw $v1,0x0008($a0)
		136: Instruct <= 32'b000000_11010_00000_00000_00000_001000;//jr $26
		*/
		
		/*
		0: Instruct <= 32'b000010_00000000000000000000000011; //j Normal
		1: Instruct <= 32'b000010_00000000000000000000011110; //j Interrupt
		2: Instruct <= 32'b000010_00000000000000000000100110; //j Exit
		3: Instruct <= 32'b001111_00000_00100_1000000000000000;  //lui $a0,0x80000000
		4: Instruct <= 32'b001111_00000_00010_0000000000000000;  //lui $v0,0
		5: Instruct <= 32'b001111_00000_00011_0000000000000000;  //lui $v0,0
		6: Instruct <= 32'b000000_00000_00000_01000_00000_100000;//add $t0,$0,$0
		7: Instruct <= 32'b000000_00000_00000_01001_00000_100000;//add $t1,$0,$0
		8: Instruct <= 32'b001000_00000_00010_0000000000000010;  //addi $v0,$0,0x0002
		9: Instruct <= 32'b001000_00000_00011_0000000000001010;  //addi $v1,$0,0x000a
		10: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		11: Instruct <= 32'b100011_00100_01000_0000000000100000;   //loop1: lw $t0,0x0020($a0)
		12: Instruct <= 32'b000100_01000_00011_0000000000000001;  //beq $t0,$v1,break1
		13: Instruct <= 32'b000010_00000000000000000000001011;    // j loop1 
		14: Instruct <= 32'b100011_00100_01001_0000000000011100;  //break1: lw $t1,0x001c($a0)
		15: Instruct <= 32'b001000_00000_00010_0000000000000000;  //addi $v0,$0,0x0
		16: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		17: Instruct <= 32'b000000_00000_01001_10000_00000_100000; //add $s0,$0,$t1
		18: Instruct <= 32'b001000_00000_00010_0000000000000010;  //addi $v0,$0,0x0002
		19: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		20: Instruct <= 32'b100011_00100_01000_0000000000100000;   //loop2: lw $t0,0x0020($a0)
		21: Instruct <= 32'b000100_01000_00011_0000000000000001;  //beq $t0,$v1,break2
		22: Instruct <= 32'b000010_00000000000000000000010100;    // j loop2 
		23: Instruct <= 32'b100011_00100_01001_0000000000011100;  //break2: lw $t1,0x001c($a0)
		24: Instruct <= 32'b001000_00000_00010_0000000000000000;  //addi $v0,$0,0x0
		25: Instruct <= 32'b101011_00100_00010_0000000000100000; //sw $v0,0x0020($a0)
		26: Instruct <= 32'b000000_00000_01001_10001_00000_100000; //add $s1,$0,$t1
		
		27: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		28: Instruct <= 32'b000100_00000_10010_0000000000000111; //compare: beq $0,$s2,result
		29: Instruct <= 32'b000001_10010_00000_0000000000000011; //bltz $s2,neg
		30: Instruct <= 32'b000000_10000_10001_10000_00000_100010; //pos: sub $s0,$s0,$s1
		31: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		32: Instruct <= 32'b000010_00000000000000000000011100;    // j compare
		33: Instruct <= 32'b000000_10001_10000_10001_00000_100010; //neg: sub $s1,$s1,$s0
		34: Instruct <= 32'b000000_10000_10001_10010_00000_100010; //sub $s2,$s0,$s1
		35: Instruct <= 32'b000010_00000000000000000000011100;    // j compare
		36: Instruct <= 32'b101011_00100_10000_0000000000011000;  // result: sw $s0,00x0018($a0)
		37: Instruct <= 32'b001000_00000_00010_0000000000000001;  //addi $v0,$0,0x0001
		38: Instruct <= 32'b001000_00000_00011_0000000000000101;  //addi $v1,$0,0x0005
		39: Instruct <= 32'b101011_00100_00010_0000000000100000;  //sw $v0,0x0020($a0)
		40: Instruct <= 32'b100011_00100_01010_0000000000100000;   //loop3: lw $t2,0x0020($a0)
		41: Instruct <= 32'b000100_01010_00011_0000000000000001;  //beq $t2,$v1,break3
		42: Instruct <= 32'b000010_00000000000000000000101000;    // j loop3
		43: Instruct <= 32'b001000_00000_00010_0000000000000000;  //break3:addi $v0,$0,0x0000
		44: Instruct <= 32'b101011_00100_00010_0000000000100000;  //sw $v0,0x0020($a0)
		45: Instruct <= 32'b001111_00000_00100_0100000000000000;  //lui $a0,0x40000000
		46: Instruct <= 32'b101011_00100_10000_0000000000001100;  //sw $s0,0x000c($a0) 
		*/
		/*
		0: Instruct <= 32'b001000_00000_00100_0000000000000001; //addi $a0, $0, 1
		1: Instruct <= 32'b0;
		2: Instruct <= 32'b001000_00000_00101_0000000000000001; //addi $a1, $0, 1
		3: Instruct <= 32'b001000_00000_00110_0000000000000010; //addi $a2, $0, 2		
		4: Instruct <= 32'b000000_00101_00100_00101_00000_100000; //add $a1, $a1, $a0
		5: Instruct <= 32'b000100_00101_00110_1111111111111110; //beq $a1, $a2, -2
		6: Instruct <= 32'b0; //nop
		*/
		/*
		// beq_test
		0: Instruct <= 32'b001000_00000_00100_0000000000000001; //addi $a0, $0, 1
		1: Instruct <= 32'b001000_00000_00101_0000000000000001;//addi $a1, $0, 1
		2: Instruct <= 32'b0; //nop
		3: Instruct <= 32'b0; //nop
		4: Instruct <= 32'b001000_00000_00110_0000000000000010; //addi $a2, $0, 2: 
		5: Instruct <= 32'b0; //nop
		6: Instruct <= 32'b000000_00101_00100_00101_00000_100000; //add $a1, $a1, $a0
		7: Instruct <= 32'b0; //nop
		8: Instruct <= 32'b0; //nop
		9: Instruct <= 32'b000100_00000_00000_1111111111111100; //beq $0, $0, -4
		10: Instruct <= 32'b000000_00101_00100_00110_00000_100000; //add $a2, $a1, $a0
		11: Instruct <= 32'b000000_00101_00100_00110_00000_100000; //add $a2, $a1, $a0
		12: Instruct <= 32'b000000_00101_00100_00110_00000_100000; //add $a2, $a1, $a0
		*/
	   default:	Instruct <= 32'h0000_0000; // nop
	endcase
	end
end
endmodule
